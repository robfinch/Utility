`timescale 1ns / 1ps
// ============================================================================
//        __
//   \\__/ o\    (C) 2013-2022  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
// BusError.v
// - generate a bus timeout error if a cycle has been active without an ack
//   for too long of a time.
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// ============================================================================
//
module BusError(rst_i, clk_i, cyc_i, ack_i, stb_i, adr_i, err_o);
parameter pTO=28'd250;
input rst_i;
input clk_i;
input cyc_i;
input ack_i;
input stb_i;
input [31:0] adr_i;
output err_o;
reg err_o;

reg [27:0] tocnt;

always_ff @(posedge clk_i)
if (rst_i) begin
	err_o <= 1'b0;
	tocnt <= 28'd1;
end
else begin
	err_o <= 1'b0;
	// If there is no bus cycle active, or if the bus cycle
	// has been acknowledged, reset the timeout count.
	if (ack_i || !cyc_i) begin
		tocnt <= 28'd1;
		err_o <= 1'b0;
	end
	else if (tocnt < pTO)
		tocnt <= tocnt + 28'd1;
	else if (cyc_i && stb_i && (adr_i[31:4]==28'hFFDCFFE)) begin	// conflist with configrec ?
		tocnt <= 28'd1;
		err_o <= 1'b0;
	end
	else
		err_o <= 1'b1;
end

endmodule
